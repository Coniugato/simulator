`timescale 1ns / 100ps

// convert unsigned integer to float
module fcvt_s_wu(
    input wire [31:0] x,
    output wire [31:0] y,
    input clk);

    wire [32:0] xs =
        x[31] ? (x[7] ? ({1'b0, x} + (33'b1<<8)) : {1'b0, x}) :
        x[30] ? (x[6] ? ({1'b0, x} + (33'b1<<7)) : {1'b0, x}) :
        x[29] ? (x[5] ? ({1'b0, x} + (33'b1<<6)) : {1'b0, x}) :
        x[28] ? (x[4] ? ({1'b0, x} + (33'b1<<5)) : {1'b0, x}) :
        x[27] ? (x[3] ? ({1'b0, x} + (33'b1<<4)) : {1'b0, x}) :
        x[26] ? (x[2] ? ({1'b0, x} + (33'b1<<3)) : {1'b0, x}) :
        x[25] ? (x[1] ? ({1'b0, x} + (33'b1<<2)) : {1'b0, x}) :
        x[24] ? (x[0] ? ({1'b0, x} + (33'b1<<1)) : {1'b0, x}) :
        {1'b0, x};

    assign y =
        xs[32] ? {1'b0, 8'd159, xs[31:9]} : 
        xs[31] ? {1'b0, 8'd158, xs[30:8]} :
        xs[30] ? {1'b0, 8'd157, xs[29:7]} :
        xs[29] ? {1'b0, 8'd156, xs[28:6]} :
        xs[28] ? {1'b0, 8'd155, xs[27:5]} :
        xs[27] ? {1'b0, 8'd154, xs[26:4]} :
        xs[26] ? {1'b0, 8'd153, xs[25:3]} :
        xs[25] ? {1'b0, 8'd152, xs[24:2]} :
        xs[24] ? {1'b0, 8'd151, xs[23:1]} :
        xs[23] ? {1'b0, 8'd150, xs[22:0]} :
        xs[22] ? {1'b0, 8'd149, xs[21:0], 1'b0} :
        xs[21] ? {1'b0, 8'd148, xs[20:0], 2'b0} :
        xs[20] ? {1'b0, 8'd147, xs[19:0], 3'b0} :
        xs[19] ? {1'b0, 8'd146, xs[18:0], 4'b0} :
        xs[18] ? {1'b0, 8'd145, xs[17:0], 5'b0} :
        xs[17] ? {1'b0, 8'd144, xs[16:0], 6'b0} :
        xs[16] ? {1'b0, 8'd143, xs[15:0], 7'b0} :
        xs[15] ? {1'b0, 8'd142, xs[14:0], 8'b0} :
        xs[14] ? {1'b0, 8'd141, xs[13:0], 9'b0} :
        xs[13] ? {1'b0, 8'd140, xs[12:0], 10'b0} :
        xs[12] ? {1'b0, 8'd139, xs[11:0], 11'b0} :
        xs[11] ? {1'b0, 8'd138, xs[10:0], 12'b0} :
        xs[10] ? {1'b0, 8'd137, xs[9:0], 13'b0} :
        xs[9] ? {1'b0, 8'd136, xs[8:0], 14'b0} :
        xs[8] ? {1'b0, 8'd135, xs[7:0], 15'b0} :
        xs[7] ? {1'b0, 8'd134, xs[6:0], 16'b0} :
        xs[6] ? {1'b0, 8'd133, xs[5:0], 17'b0} :
        xs[5] ? {1'b0, 8'd132, xs[4:0], 18'b0} :
        xs[4] ? {1'b0, 8'd131, xs[3:0], 19'b0} :
        xs[3] ? {1'b0, 8'd130, xs[2:0], 20'b0} :
        xs[2] ? {1'b0, 8'd129, xs[1:0], 21'b0} :
        xs[1] ? {1'b0, 8'd128, xs[0], 22'b0} :
        xs[0] ? {1'b0, 8'd127, 23'b0} :
        32'b0;
endmodule